library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity seno is
  port (
    ADDR : in  std_logic_vector(7 downto 0);
    CLK  : in  std_logic;
    DOUT : out std_logic_vector(7 downto 0) );
end seno;

architecture rtl of seno is
 
  type cell is array (0 to 255) of std_logic_vector(7 downto 0);
  constant memoria  : cell := (
  0  => x"00", 
 1  => x"00", 
 2  => x"00", 
 3  => x"00", 
 4  => x"00", 
 5  => x"00", 
 6  => x"01", 
 7  => x"01", 
 8  => x"02", 
 9  => x"03", 
 10  => x"03", 
 11  => x"04", 
 12  => x"05", 
 13  => x"06", 
 14  => x"07", 
 15  => x"08", 
 16  => x"09", 
 17  => x"0B", 
 18  => x"0C", 
 19  => x"0D", 
 20  => x"0F", 
 21  => x"10", 
 22  => x"12", 
 23  => x"13", 
 24  => x"15", 
 25  => x"17", 
 26  => x"19", 
 27  => x"1B", 
 28  => x"1D", 
 29  => x"1F", 
 30  => x"21", 
 31  => x"23", 
 32  => x"25", 
 33  => x"27", 
 34  => x"2A", 
 35  => x"2C", 
 36  => x"2E", 
 37  => x"31", 
 38  => x"33", 
 39  => x"36", 
 40  => x"39", 
 41  => x"3B", 
 42  => x"3E", 
 43  => x"41", 
 44  => x"43", 
 45  => x"46", 
 46  => x"49", 
 47  => x"4C", 
 48  => x"4F", 
 49  => x"52", 
 50  => x"55", 
 51  => x"58", 
 52  => x"5B", 
 53  => x"5E", 
 54  => x"61", 
 55  => x"64", 
 56  => x"67", 
 57  => x"6A", 
 58  => x"6D", 
 59  => x"70", 
 60  => x"73", 
 61  => x"76", 
 62  => x"7A", 
 63  => x"7D", 
 64  => x"80", 
 65  => x"83", 
 66  => x"86", 
 67  => x"89", 
 68  => x"8C", 
 69  => x"8F", 
 70  => x"93", 
 71  => x"96", 
 72  => x"99", 
 73  => x"9C", 
 74  => x"9F", 
 75  => x"A2", 
 76  => x"A5", 
 77  => x"A8", 
 78  => x"AB", 
 79  => x"AE", 
 80  => x"B1", 
 81  => x"B4", 
 82  => x"B6", 
 83  => x"B9", 
 84  => x"BC", 
 85  => x"BF", 
 86  => x"C1", 
 87  => x"C4", 
 88  => x"C7", 
 89  => x"C9", 
 90  => x"CC", 
 91  => x"CE", 
 92  => x"D1", 
 93  => x"D3", 
 94  => x"D5", 
 95  => x"D8", 
 96  => x"DA", 
 97  => x"DC", 
 98  => x"DE", 
 99  => x"E0", 
 100  => x"E2", 
 101  => x"E4", 
 102  => x"E6", 
 103  => x"E8", 
 104  => x"EA", 
 105  => x"EB", 
 106  => x"ED", 
 107  => x"EF", 
 108  => x"F0", 
 109  => x"F1", 
 110  => x"F3", 
 111  => x"F4", 
 112  => x"F5", 
 113  => x"F6", 
 114  => x"F8", 
 115  => x"F9", 
 116  => x"F9", 
 117  => x"FA", 
 118  => x"FB", 
 119  => x"FC", 
 120  => x"FC", 
 121  => x"FD", 
 122  => x"FD", 
 123  => x"FE", 
 124  => x"FE", 
 125  => x"FE", 
 126  => x"FE", 
 127  => x"FE", 
 128  => x"FE", 
 129  => x"FE", 
 130  => x"FE", 
 131  => x"FE", 
 132  => x"FE", 
 133  => x"FD", 
 134  => x"FD", 
 135  => x"FC", 
 136  => x"FC", 
 137  => x"FB", 
 138  => x"FA", 
 139  => x"F9", 
 140  => x"F9", 
 141  => x"F8", 
 142  => x"F6", 
 143  => x"F5", 
 144  => x"F4", 
 145  => x"F3", 
 146  => x"F1", 
 147  => x"F0", 
 148  => x"EF", 
 149  => x"ED", 
 150  => x"EB", 
 151  => x"EA", 
 152  => x"E8", 
 153  => x"E6", 
 154  => x"E4", 
 155  => x"E2", 
 156  => x"E0", 
 157  => x"DE", 
 158  => x"DC", 
 159  => x"DA", 
 160  => x"D8", 
 161  => x"D5", 
 162  => x"D3", 
 163  => x"D1", 
 164  => x"CE", 
 165  => x"CC", 
 166  => x"C9", 
 167  => x"C7", 
 168  => x"C4", 
 169  => x"C1", 
 170  => x"BF", 
 171  => x"BC", 
 172  => x"B9", 
 173  => x"B6", 
 174  => x"B4", 
 175  => x"B1", 
 176  => x"AE", 
 177  => x"AB", 
 178  => x"A8", 
 179  => x"A5", 
 180  => x"A2", 
 181  => x"9F", 
 182  => x"9C", 
 183  => x"99", 
 184  => x"96", 
 185  => x"93", 
 186  => x"8F", 
 187  => x"8C", 
 188  => x"89", 
 189  => x"86", 
 190  => x"83", 
 191  => x"80", 
 192  => x"7D", 
 193  => x"7A", 
 194  => x"76", 
 195  => x"73", 
 196  => x"70", 
 197  => x"6D", 
 198  => x"6A", 
 199  => x"67", 
 200  => x"64", 
 201  => x"61", 
 202  => x"5E", 
 203  => x"5B", 
 204  => x"58", 
 205  => x"55", 
 206  => x"52", 
 207  => x"4F", 
 208  => x"4C", 
 209  => x"49", 
 210  => x"46", 
 211  => x"43", 
 212  => x"41", 
 213  => x"3E", 
 214  => x"3B", 
 215  => x"39", 
 216  => x"36", 
 217  => x"33", 
 218  => x"31", 
 219  => x"2E", 
 220  => x"2C", 
 221  => x"2A", 
 222  => x"27", 
 223  => x"25", 
 224  => x"23", 
 225  => x"21", 
 226  => x"1F", 
 227  => x"1D", 
 228  => x"1B", 
 229  => x"19", 
 230  => x"17", 
 231  => x"15", 
 232  => x"13", 
 233  => x"12", 
 234  => x"10", 
 235  => x"0F", 
 236  => x"0D", 
 237  => x"0C", 
 238  => x"0B", 
 239  => x"09", 
 240  => x"08", 
 241  => x"07", 
 242  => x"06", 
 243  => x"05", 
 244  => x"04", 
 245  => x"03", 
 246  => x"03", 
 247  => x"02", 
 248  => x"01", 
 249  => x"01", 
 250  => x"00", 
 251  => x"00", 
 252  => x"00", 
 253  => x"00", 
 254  => x"00", 
 255  => x"00"); 

  
begin
  
  process (clk)
  begin 
    if clk'event and clk = '1' then 
      DOUT<=memoria(to_integer(unsigned(addr)));
    end if;
  end process;
 
end rtl;
